// Video_System.v

// Generated using ACDS version 14.0 200 at 2015.05.06.01:36:28

`timescale 1 ps / 1 ps
module Video_System (
		inout  wire [15:0] SRAM_DQ_to_and_from_the_Pixel_Buffer, //   Pixel_Buffer_external_interface.DQ
		output wire [19:0] SRAM_ADDR_from_the_Pixel_Buffer,      //                                  .ADDR
		output wire        SRAM_LB_N_from_the_Pixel_Buffer,      //                                  .LB_N
		output wire        SRAM_UB_N_from_the_Pixel_Buffer,      //                                  .UB_N
		output wire        SRAM_CE_N_from_the_Pixel_Buffer,      //                                  .CE_N
		output wire        SRAM_OE_N_from_the_Pixel_Buffer,      //                                  .OE_N
		output wire        SRAM_WE_N_from_the_Pixel_Buffer,      //                                  .WE_N
		output wire        VGA_CLK_from_the_VGA_Controller,      // VGA_Controller_external_interface.CLK
		output wire        VGA_HS_from_the_VGA_Controller,       //                                  .HS
		output wire        VGA_VS_from_the_VGA_Controller,       //                                  .VS
		output wire        VGA_BLANK_from_the_VGA_Controller,    //                                  .BLANK
		output wire        VGA_SYNC_from_the_VGA_Controller,     //                                  .SYNC
		output wire [7:0]  VGA_R_from_the_VGA_Controller,        //                                  .R
		output wire [7:0]  VGA_G_from_the_VGA_Controller,        //                                  .G
		output wire [7:0]  VGA_B_from_the_VGA_Controller,        //                                  .B
		input  wire        clk_0,                                //                      clk_0_clk_in.clk
		input  wire        reset_n,                              //                clk_0_clk_in_reset.reset_n
		input  wire [7:0]  keycode_export,                       //                           keycode.export
		output wire        sdram_out_clk_clk,                    //                     sdram_out_clk.clk
		output wire [12:0] sdram_wire_addr,                      //                        sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                        //                                  .ba
		output wire        sdram_wire_cas_n,                     //                                  .cas_n
		output wire        sdram_wire_cke,                       //                                  .cke
		output wire        sdram_wire_cs_n,                      //                                  .cs_n
		inout  wire [31:0] sdram_wire_dq,                        //                                  .dq
		output wire [3:0]  sdram_wire_dqm,                       //                                  .dqm
		output wire        sdram_wire_ras_n,                     //                                  .ras_n
		output wire        sdram_wire_we_n,                      //                                  .we_n
		input  wire [7:0]  press_export                          //                             press.export
	);

	wire         alpha_blender_avalon_blended_source_endofpacket;                             // Alpha_Blender:output_endofpacket -> Dual_Clock_FIFO:stream_in_endofpacket
	wire         alpha_blender_avalon_blended_source_valid;                                   // Alpha_Blender:output_valid -> Dual_Clock_FIFO:stream_in_valid
	wire         alpha_blender_avalon_blended_source_startofpacket;                           // Alpha_Blender:output_startofpacket -> Dual_Clock_FIFO:stream_in_startofpacket
	wire  [29:0] alpha_blender_avalon_blended_source_data;                                    // Alpha_Blender:output_data -> Dual_Clock_FIFO:stream_in_data
	wire         alpha_blender_avalon_blended_source_ready;                                   // Dual_Clock_FIFO:stream_in_ready -> Alpha_Blender:output_ready
	wire         char_buffer_with_dma_avalon_char_source_endofpacket;                         // Char_Buffer_with_DMA:stream_endofpacket -> Alpha_Blender:foreground_endofpacket
	wire         char_buffer_with_dma_avalon_char_source_valid;                               // Char_Buffer_with_DMA:stream_valid -> Alpha_Blender:foreground_valid
	wire         char_buffer_with_dma_avalon_char_source_startofpacket;                       // Char_Buffer_with_DMA:stream_startofpacket -> Alpha_Blender:foreground_startofpacket
	wire  [39:0] char_buffer_with_dma_avalon_char_source_data;                                // Char_Buffer_with_DMA:stream_data -> Alpha_Blender:foreground_data
	wire         char_buffer_with_dma_avalon_char_source_ready;                               // Alpha_Blender:foreground_ready -> Char_Buffer_with_DMA:stream_ready
	wire         dual_clock_fifo_avalon_dc_buffer_source_endofpacket;                         // Dual_Clock_FIFO:stream_out_endofpacket -> VGA_Controller:endofpacket
	wire         dual_clock_fifo_avalon_dc_buffer_source_valid;                               // Dual_Clock_FIFO:stream_out_valid -> VGA_Controller:valid
	wire         dual_clock_fifo_avalon_dc_buffer_source_startofpacket;                       // Dual_Clock_FIFO:stream_out_startofpacket -> VGA_Controller:startofpacket
	wire  [29:0] dual_clock_fifo_avalon_dc_buffer_source_data;                                // Dual_Clock_FIFO:stream_out_data -> VGA_Controller:data
	wire         dual_clock_fifo_avalon_dc_buffer_source_ready;                               // VGA_Controller:ready -> Dual_Clock_FIFO:stream_out_ready
	wire         pixel_buffer_dma_avalon_pixel_source_endofpacket;                            // Pixel_Buffer_DMA:stream_endofpacket -> Pixel_RGB_Resampler:stream_in_endofpacket
	wire         pixel_buffer_dma_avalon_pixel_source_valid;                                  // Pixel_Buffer_DMA:stream_valid -> Pixel_RGB_Resampler:stream_in_valid
	wire         pixel_buffer_dma_avalon_pixel_source_startofpacket;                          // Pixel_Buffer_DMA:stream_startofpacket -> Pixel_RGB_Resampler:stream_in_startofpacket
	wire  [15:0] pixel_buffer_dma_avalon_pixel_source_data;                                   // Pixel_Buffer_DMA:stream_data -> Pixel_RGB_Resampler:stream_in_data
	wire         pixel_buffer_dma_avalon_pixel_source_ready;                                  // Pixel_RGB_Resampler:stream_in_ready -> Pixel_Buffer_DMA:stream_ready
	wire         pixel_rgb_resampler_avalon_rgb_source_endofpacket;                           // Pixel_RGB_Resampler:stream_out_endofpacket -> Pixel_Scaler:stream_in_endofpacket
	wire         pixel_rgb_resampler_avalon_rgb_source_valid;                                 // Pixel_RGB_Resampler:stream_out_valid -> Pixel_Scaler:stream_in_valid
	wire         pixel_rgb_resampler_avalon_rgb_source_startofpacket;                         // Pixel_RGB_Resampler:stream_out_startofpacket -> Pixel_Scaler:stream_in_startofpacket
	wire  [29:0] pixel_rgb_resampler_avalon_rgb_source_data;                                  // Pixel_RGB_Resampler:stream_out_data -> Pixel_Scaler:stream_in_data
	wire         pixel_rgb_resampler_avalon_rgb_source_ready;                                 // Pixel_Scaler:stream_in_ready -> Pixel_RGB_Resampler:stream_out_ready
	wire         pixel_scaler_avalon_scaler_source_endofpacket;                               // Pixel_Scaler:stream_out_endofpacket -> Alpha_Blender:background_endofpacket
	wire         pixel_scaler_avalon_scaler_source_valid;                                     // Pixel_Scaler:stream_out_valid -> Alpha_Blender:background_valid
	wire         pixel_scaler_avalon_scaler_source_startofpacket;                             // Pixel_Scaler:stream_out_startofpacket -> Alpha_Blender:background_startofpacket
	wire  [29:0] pixel_scaler_avalon_scaler_source_data;                                      // Pixel_Scaler:stream_out_data -> Alpha_Blender:background_data
	wire         pixel_scaler_avalon_scaler_source_ready;                                     // Alpha_Blender:background_ready -> Pixel_Scaler:stream_out_ready
	wire         video_pll_0_vga_clk_clk;                                                     // video_pll_0:vga_clk_clk -> [Dual_Clock_FIFO:clk_stream_out, VGA_Controller:clk, rst_controller_002:clk, rst_controller_003:clk]
	wire         cpu_data_master_waitrequest;                                                 // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                                   // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [28:0] cpu_data_master_address;                                                     // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire         cpu_data_master_write;                                                       // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire         cpu_data_master_read;                                                        // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                                    // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_debugaccess;                                                 // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                                  // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_instruction_master_waitrequest;                                          // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [28:0] cpu_instruction_master_address;                                              // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                                 // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                             // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         pixel_buffer_dma_avalon_pixel_dma_master_waitrequest;                        // mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_waitrequest -> Pixel_Buffer_DMA:master_waitrequest
	wire  [31:0] pixel_buffer_dma_avalon_pixel_dma_master_address;                            // Pixel_Buffer_DMA:master_address -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_address
	wire         pixel_buffer_dma_avalon_pixel_dma_master_lock;                               // Pixel_Buffer_DMA:master_arbiterlock -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_lock
	wire         pixel_buffer_dma_avalon_pixel_dma_master_read;                               // Pixel_Buffer_DMA:master_read -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_read
	wire  [15:0] pixel_buffer_dma_avalon_pixel_dma_master_readdata;                           // mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_readdata -> Pixel_Buffer_DMA:master_readdata
	wire         pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid;                      // mm_interconnect_0:Pixel_Buffer_DMA_avalon_pixel_dma_master_readdatavalid -> Pixel_Buffer_DMA:master_readdatavalid
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_waitrequest; // Char_Buffer_with_DMA:buf_waitrequest -> mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_waitrequest
	wire   [7:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_writedata -> Char_Buffer_with_DMA:buf_writedata
	wire  [12:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_address;     // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_address -> Char_Buffer_with_DMA:buf_address
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_chipselect -> Char_Buffer_with_DMA:buf_chipselect
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_write;       // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_write -> Char_Buffer_with_DMA:buf_write
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_read;        // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_read -> Char_Buffer_with_DMA:buf_read
	wire   [7:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_readdata;    // Char_Buffer_with_DMA:buf_readdata -> mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_readdata
	wire   [0:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_buffer_slave_byteenable -> Char_Buffer_with_DMA:buf_byteenable
	wire  [31:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_writedata;  // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_writedata -> Char_Buffer_with_DMA:ctrl_writedata
	wire   [0:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_address;    // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_address -> Char_Buffer_with_DMA:ctrl_address
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_chipselect; // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_chipselect -> Char_Buffer_with_DMA:ctrl_chipselect
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_write;      // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_write -> Char_Buffer_with_DMA:ctrl_write
	wire         mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_read;       // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_read -> Char_Buffer_with_DMA:ctrl_read
	wire  [31:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_readdata;   // Char_Buffer_with_DMA:ctrl_readdata -> mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_readdata
	wire   [3:0] mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_byteenable; // mm_interconnect_0:Char_Buffer_with_DMA_avalon_char_control_slave_byteenable -> Char_Buffer_with_DMA:ctrl_byteenable
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata;           // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_writedata -> Pixel_Buffer_DMA:slave_writedata
	wire   [1:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address;             // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_address -> Pixel_Buffer_DMA:slave_address
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write;               // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_write -> Pixel_Buffer_DMA:slave_write
	wire         mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read;                // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_read -> Pixel_Buffer_DMA:slave_read
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata;            // Pixel_Buffer_DMA:slave_readdata -> mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_readdata
	wire   [3:0] mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable;          // mm_interconnect_0:Pixel_Buffer_DMA_avalon_control_slave_byteenable -> Pixel_Buffer_DMA:slave_byteenable
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata;                  // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_writedata -> Pixel_Buffer:writedata
	wire  [19:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_address;                    // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_address -> Pixel_Buffer:address
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_write;                      // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_write -> Pixel_Buffer:write
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_read;                       // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_read -> Pixel_Buffer:read
	wire  [15:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata;                   // Pixel_Buffer:readdata -> mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_readdata
	wire         mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid;              // Pixel_Buffer:readdatavalid -> mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_readdatavalid
	wire   [1:0] mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable;                 // mm_interconnect_0:Pixel_Buffer_avalon_sram_slave_byteenable -> Pixel_Buffer:byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                         // CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                           // mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                             // mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                               // mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                                // mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                            // CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                         // mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                          // mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire   [1:0] mm_interconnect_0_keycode_s1_address;                                        // mm_interconnect_0:keycode_s1_address -> keycode:address
	wire  [31:0] mm_interconnect_0_keycode_s1_readdata;                                       // keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	wire  [31:0] mm_interconnect_0_sdram_clk_pll_slave_writedata;                             // mm_interconnect_0:sdram_clk_pll_slave_writedata -> sdram_clk:writedata
	wire   [1:0] mm_interconnect_0_sdram_clk_pll_slave_address;                               // mm_interconnect_0:sdram_clk_pll_slave_address -> sdram_clk:address
	wire         mm_interconnect_0_sdram_clk_pll_slave_write;                                 // mm_interconnect_0:sdram_clk_pll_slave_write -> sdram_clk:write
	wire         mm_interconnect_0_sdram_clk_pll_slave_read;                                  // mm_interconnect_0:sdram_clk_pll_slave_read -> sdram_clk:read
	wire  [31:0] mm_interconnect_0_sdram_clk_pll_slave_readdata;                              // sdram_clk:readdata -> mm_interconnect_0:sdram_clk_pll_slave_readdata
	wire         mm_interconnect_0_sdram_controller_0_s1_waitrequest;                         // sdram_controller_0:za_waitrequest -> mm_interconnect_0:sdram_controller_0_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_controller_0_s1_writedata;                           // mm_interconnect_0:sdram_controller_0_s1_writedata -> sdram_controller_0:az_data
	wire  [24:0] mm_interconnect_0_sdram_controller_0_s1_address;                             // mm_interconnect_0:sdram_controller_0_s1_address -> sdram_controller_0:az_addr
	wire         mm_interconnect_0_sdram_controller_0_s1_chipselect;                          // mm_interconnect_0:sdram_controller_0_s1_chipselect -> sdram_controller_0:az_cs
	wire         mm_interconnect_0_sdram_controller_0_s1_write;                               // mm_interconnect_0:sdram_controller_0_s1_write -> sdram_controller_0:az_wr_n
	wire         mm_interconnect_0_sdram_controller_0_s1_read;                                // mm_interconnect_0:sdram_controller_0_s1_read -> sdram_controller_0:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_controller_0_s1_readdata;                            // sdram_controller_0:za_data -> mm_interconnect_0:sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_sdram_controller_0_s1_readdatavalid;                       // sdram_controller_0:za_valid -> mm_interconnect_0:sdram_controller_0_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_controller_0_s1_byteenable;                          // mm_interconnect_0:sdram_controller_0_s1_byteenable -> sdram_controller_0:az_be_n
	wire   [1:0] mm_interconnect_0_press_s1_address;                                          // mm_interconnect_0:press_s1_address -> press:address
	wire  [31:0] mm_interconnect_0_press_s1_readdata;                                         // press:readdata -> mm_interconnect_0:press_s1_readdata
	wire  [31:0] cpu_d_irq_irq;                                                               // irq_mapper:sender_irq -> CPU:d_irq
	wire         rst_controller_reset_out_reset;                                              // rst_controller:reset_out -> [Alpha_Blender:reset, Char_Buffer_with_DMA:reset, Pixel_Buffer:reset, Pixel_Buffer_DMA:reset, Pixel_RGB_Resampler:reset, Pixel_Scaler:reset, mm_interconnect_0:Pixel_Buffer_DMA_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                          // rst_controller_001:reset_out -> [CPU:reset_n, Dual_Clock_FIFO:reset_stream_in, irq_mapper:reset, keycode:reset_n, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, press:reset_n, rst_translator:in_reset, sdram_clk:reset, video_pll_0:ref_reset_reset]
	wire         rst_controller_001_reset_out_reset_req;                                      // rst_controller_001:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                           // CPU:jtag_debug_module_resetrequest -> [rst_controller_001:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in0]
	wire         rst_controller_002_reset_out_reset;                                          // rst_controller_002:reset_out -> Dual_Clock_FIFO:reset_stream_out
	wire         video_pll_0_reset_source_reset;                                              // video_pll_0:reset_source_reset -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	wire         rst_controller_003_reset_out_reset;                                          // rst_controller_003:reset_out -> VGA_Controller:reset
	wire         rst_controller_004_reset_out_reset;                                          // rst_controller_004:reset_out -> [mm_interconnect_0:sdram_controller_0_reset_reset_bridge_in_reset_reset, sdram_controller_0:reset_n]

	Video_System_Alpha_Blender alpha_blender (
		.clk                      (clk_0),                                                 //                    clk.clk
		.reset                    (rst_controller_reset_out_reset),                        //                  reset.reset
		.foreground_data          (char_buffer_with_dma_avalon_char_source_data),          // avalon_foreground_sink.data
		.foreground_startofpacket (char_buffer_with_dma_avalon_char_source_startofpacket), //                       .startofpacket
		.foreground_endofpacket   (char_buffer_with_dma_avalon_char_source_endofpacket),   //                       .endofpacket
		.foreground_valid         (char_buffer_with_dma_avalon_char_source_valid),         //                       .valid
		.foreground_ready         (char_buffer_with_dma_avalon_char_source_ready),         //                       .ready
		.background_data          (pixel_scaler_avalon_scaler_source_data),                // avalon_background_sink.data
		.background_startofpacket (pixel_scaler_avalon_scaler_source_startofpacket),       //                       .startofpacket
		.background_endofpacket   (pixel_scaler_avalon_scaler_source_endofpacket),         //                       .endofpacket
		.background_valid         (pixel_scaler_avalon_scaler_source_valid),               //                       .valid
		.background_ready         (pixel_scaler_avalon_scaler_source_ready),               //                       .ready
		.output_ready             (alpha_blender_avalon_blended_source_ready),             //  avalon_blended_source.ready
		.output_data              (alpha_blender_avalon_blended_source_data),              //                       .data
		.output_startofpacket     (alpha_blender_avalon_blended_source_startofpacket),     //                       .startofpacket
		.output_endofpacket       (alpha_blender_avalon_blended_source_endofpacket),       //                       .endofpacket
		.output_valid             (alpha_blender_avalon_blended_source_valid)              //                       .valid
	);

	Video_System_CPU cpu (
		.clk                                   (clk_0),                                               //                       clk.clk
		.reset_n                               (~rst_controller_001_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_001_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	Video_System_Char_Buffer_with_DMA char_buffer_with_dma (
		.clk                  (clk_0),                                                                       //                       clk.clk
		.reset                (rst_controller_reset_out_reset),                                              //                     reset.reset
		.ctrl_address         (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (char_buffer_with_dma_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (char_buffer_with_dma_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (char_buffer_with_dma_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (char_buffer_with_dma_avalon_char_source_valid),                               //                          .valid
		.stream_data          (char_buffer_with_dma_avalon_char_source_data)                                 //                          .data
	);

	Video_System_Dual_Clock_FIFO dual_clock_fifo (
		.clk_stream_in            (clk_0),                                                 //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_001_reset_out_reset),                    //         reset_stream_in.reset
		.clk_stream_out           (video_pll_0_vga_clk_clk),                               //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                    //        reset_stream_out.reset
		.stream_in_ready          (alpha_blender_avalon_blended_source_ready),             //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blender_avalon_blended_source_startofpacket),     //                        .startofpacket
		.stream_in_endofpacket    (alpha_blender_avalon_blended_source_endofpacket),       //                        .endofpacket
		.stream_in_valid          (alpha_blender_avalon_blended_source_valid),             //                        .valid
		.stream_in_data           (alpha_blender_avalon_blended_source_data),              //                        .data
		.stream_out_ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (dual_clock_fifo_avalon_dc_buffer_source_data)           //                        .data
	);

	Video_System_Pixel_Buffer pixel_buffer (
		.clk           (clk_0),                                                          //                clk.clk
		.reset         (rst_controller_reset_out_reset),                                 //              reset.reset
		.SRAM_DQ       (SRAM_DQ_to_and_from_the_Pixel_Buffer),                           // external_interface.export
		.SRAM_ADDR     (SRAM_ADDR_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_LB_N     (SRAM_LB_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_UB_N     (SRAM_UB_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_CE_N     (SRAM_CE_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_OE_N     (SRAM_OE_N_from_the_Pixel_Buffer),                                //                   .export
		.SRAM_WE_N     (SRAM_WE_N_from_the_Pixel_Buffer),                                //                   .export
		.address       (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	Video_System_Pixel_Buffer_DMA pixel_buffer_dma (
		.clk                  (clk_0),                                                              //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                     //                   reset.reset
		.master_readdatavalid (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_dma_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_dma_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_dma_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_dma_avalon_pixel_source_data)                           //                        .data
	);

	Video_System_Pixel_RGB_Resampler pixel_rgb_resampler (
		.clk                      (clk_0),                                               //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_avalon_pixel_source_startofpacket),  //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_avalon_pixel_source_endofpacket),    //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_avalon_pixel_source_valid),          //                  .valid
		.stream_in_ready          (pixel_buffer_dma_avalon_pixel_source_ready),          //                  .ready
		.stream_in_data           (pixel_buffer_dma_avalon_pixel_source_data),           //                  .data
		.stream_out_ready         (pixel_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (pixel_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (pixel_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (pixel_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	Video_System_Pixel_Scaler pixel_scaler (
		.clk                      (clk_0),                                               //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                reset.reset
		.stream_in_startofpacket  (pixel_rgb_resampler_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (pixel_rgb_resampler_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (pixel_rgb_resampler_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (pixel_rgb_resampler_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (pixel_rgb_resampler_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (pixel_scaler_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (pixel_scaler_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (pixel_scaler_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (pixel_scaler_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (pixel_scaler_avalon_scaler_source_data)               //                     .data
	);

	Video_System_VGA_Controller vga_controller (
		.clk           (video_pll_0_vga_clk_clk),                               //                clk.clk
		.reset         (rst_controller_003_reset_out_reset),                    //              reset.reset
		.data          (dual_clock_fifo_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (dual_clock_fifo_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (dual_clock_fifo_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (dual_clock_fifo_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (dual_clock_fifo_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (VGA_CLK_from_the_VGA_Controller),                       // external_interface.export
		.VGA_HS        (VGA_HS_from_the_VGA_Controller),                        //                   .export
		.VGA_VS        (VGA_VS_from_the_VGA_Controller),                        //                   .export
		.VGA_BLANK     (VGA_BLANK_from_the_VGA_Controller),                     //                   .export
		.VGA_SYNC      (VGA_SYNC_from_the_VGA_Controller),                      //                   .export
		.VGA_R         (VGA_R_from_the_VGA_Controller),                         //                   .export
		.VGA_G         (VGA_G_from_the_VGA_Controller),                         //                   .export
		.VGA_B         (VGA_B_from_the_VGA_Controller)                          //                   .export
	);

	Video_System_video_pll_0 video_pll_0 (
		.ref_clk_clk        (clk_0),                              //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.vga_clk_clk        (video_pll_0_vga_clk_clk),            //      vga_clk.clk
		.reset_source_reset (video_pll_0_reset_source_reset)      // reset_source.reset
	);

	Video_System_keycode keycode (
		.clk      (clk_0),                                 //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address  (mm_interconnect_0_keycode_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_keycode_s1_readdata), //                    .readdata
		.in_port  (keycode_export)                         // external_connection.export
	);

	Video_System_sdram_controller_0 sdram_controller_0 (
		.clk            (sdram_out_clk_clk),                                     //   clk.clk
		.reset_n        (~rst_controller_004_reset_out_reset),                   // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	Video_System_sdram_clk sdram_clk (
		.clk       (clk_0),                                           //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sdram_clk_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sdram_clk_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sdram_clk_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sdram_clk_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sdram_clk_pll_slave_writedata), //                      .writedata
		.c0        (sdram_out_clk_clk),                               //                    c0.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	Video_System_keycode press (
		.clk      (clk_0),                               //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_press_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_press_s1_readdata), //                    .readdata
		.in_port  (press_export)                         // external_connection.export
	);

	Video_System_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                             (clk_0),                                                                       //                                      clk_0_clk.clk
		.sdram_clk_c0_clk                                          (sdram_out_clk_clk),                                                           //                                   sdram_clk_c0.clk
		.CPU_reset_n_reset_bridge_in_reset_reset                   (rst_controller_001_reset_out_reset),                                          //              CPU_reset_n_reset_bridge_in_reset.reset
		.Pixel_Buffer_DMA_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                              //   Pixel_Buffer_DMA_reset_reset_bridge_in_reset.reset
		.sdram_controller_0_reset_reset_bridge_in_reset_reset      (rst_controller_004_reset_out_reset),                                          // sdram_controller_0_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                                   (cpu_data_master_address),                                                     //                                CPU_data_master.address
		.CPU_data_master_waitrequest                               (cpu_data_master_waitrequest),                                                 //                                               .waitrequest
		.CPU_data_master_byteenable                                (cpu_data_master_byteenable),                                                  //                                               .byteenable
		.CPU_data_master_read                                      (cpu_data_master_read),                                                        //                                               .read
		.CPU_data_master_readdata                                  (cpu_data_master_readdata),                                                    //                                               .readdata
		.CPU_data_master_write                                     (cpu_data_master_write),                                                       //                                               .write
		.CPU_data_master_writedata                                 (cpu_data_master_writedata),                                                   //                                               .writedata
		.CPU_data_master_debugaccess                               (cpu_data_master_debugaccess),                                                 //                                               .debugaccess
		.CPU_instruction_master_address                            (cpu_instruction_master_address),                                              //                         CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                        (cpu_instruction_master_waitrequest),                                          //                                               .waitrequest
		.CPU_instruction_master_read                               (cpu_instruction_master_read),                                                 //                                               .read
		.CPU_instruction_master_readdata                           (cpu_instruction_master_readdata),                                             //                                               .readdata
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_address          (pixel_buffer_dma_avalon_pixel_dma_master_address),                            //       Pixel_Buffer_DMA_avalon_pixel_dma_master.address
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_waitrequest      (pixel_buffer_dma_avalon_pixel_dma_master_waitrequest),                        //                                               .waitrequest
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_read             (pixel_buffer_dma_avalon_pixel_dma_master_read),                               //                                               .read
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_readdata         (pixel_buffer_dma_avalon_pixel_dma_master_readdata),                           //                                               .readdata
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_readdatavalid    (pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid),                      //                                               .readdatavalid
		.Pixel_Buffer_DMA_avalon_pixel_dma_master_lock             (pixel_buffer_dma_avalon_pixel_dma_master_lock),                               //                                               .lock
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_address     (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_address),     //  Char_Buffer_with_DMA_avalon_char_buffer_slave.address
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_write       (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_write),       //                                               .write
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_read        (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_read),        //                                               .read
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_readdata    (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_readdata),    //                                               .readdata
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_writedata   (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_writedata),   //                                               .writedata
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_byteenable),  //                                               .byteenable
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_waitrequest), //                                               .waitrequest
		.Char_Buffer_with_DMA_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_char_buffer_with_dma_avalon_char_buffer_slave_chipselect),  //                                               .chipselect
		.Char_Buffer_with_DMA_avalon_char_control_slave_address    (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_address),    // Char_Buffer_with_DMA_avalon_char_control_slave.address
		.Char_Buffer_with_DMA_avalon_char_control_slave_write      (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_write),      //                                               .write
		.Char_Buffer_with_DMA_avalon_char_control_slave_read       (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_read),       //                                               .read
		.Char_Buffer_with_DMA_avalon_char_control_slave_readdata   (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_readdata),   //                                               .readdata
		.Char_Buffer_with_DMA_avalon_char_control_slave_writedata  (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_writedata),  //                                               .writedata
		.Char_Buffer_with_DMA_avalon_char_control_slave_byteenable (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_byteenable), //                                               .byteenable
		.Char_Buffer_with_DMA_avalon_char_control_slave_chipselect (mm_interconnect_0_char_buffer_with_dma_avalon_char_control_slave_chipselect), //                                               .chipselect
		.CPU_jtag_debug_module_address                             (mm_interconnect_0_cpu_jtag_debug_module_address),                             //                          CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                               (mm_interconnect_0_cpu_jtag_debug_module_write),                               //                                               .write
		.CPU_jtag_debug_module_read                                (mm_interconnect_0_cpu_jtag_debug_module_read),                                //                                               .read
		.CPU_jtag_debug_module_readdata                            (mm_interconnect_0_cpu_jtag_debug_module_readdata),                            //                                               .readdata
		.CPU_jtag_debug_module_writedata                           (mm_interconnect_0_cpu_jtag_debug_module_writedata),                           //                                               .writedata
		.CPU_jtag_debug_module_byteenable                          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                          //                                               .byteenable
		.CPU_jtag_debug_module_waitrequest                         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                         //                                               .waitrequest
		.CPU_jtag_debug_module_debugaccess                         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                         //                                               .debugaccess
		.keycode_s1_address                                        (mm_interconnect_0_keycode_s1_address),                                        //                                     keycode_s1.address
		.keycode_s1_readdata                                       (mm_interconnect_0_keycode_s1_readdata),                                       //                                               .readdata
		.Pixel_Buffer_avalon_sram_slave_address                    (mm_interconnect_0_pixel_buffer_avalon_sram_slave_address),                    //                 Pixel_Buffer_avalon_sram_slave.address
		.Pixel_Buffer_avalon_sram_slave_write                      (mm_interconnect_0_pixel_buffer_avalon_sram_slave_write),                      //                                               .write
		.Pixel_Buffer_avalon_sram_slave_read                       (mm_interconnect_0_pixel_buffer_avalon_sram_slave_read),                       //                                               .read
		.Pixel_Buffer_avalon_sram_slave_readdata                   (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdata),                   //                                               .readdata
		.Pixel_Buffer_avalon_sram_slave_writedata                  (mm_interconnect_0_pixel_buffer_avalon_sram_slave_writedata),                  //                                               .writedata
		.Pixel_Buffer_avalon_sram_slave_byteenable                 (mm_interconnect_0_pixel_buffer_avalon_sram_slave_byteenable),                 //                                               .byteenable
		.Pixel_Buffer_avalon_sram_slave_readdatavalid              (mm_interconnect_0_pixel_buffer_avalon_sram_slave_readdatavalid),              //                                               .readdatavalid
		.Pixel_Buffer_DMA_avalon_control_slave_address             (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_address),             //          Pixel_Buffer_DMA_avalon_control_slave.address
		.Pixel_Buffer_DMA_avalon_control_slave_write               (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_write),               //                                               .write
		.Pixel_Buffer_DMA_avalon_control_slave_read                (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_read),                //                                               .read
		.Pixel_Buffer_DMA_avalon_control_slave_readdata            (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_readdata),            //                                               .readdata
		.Pixel_Buffer_DMA_avalon_control_slave_writedata           (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_writedata),           //                                               .writedata
		.Pixel_Buffer_DMA_avalon_control_slave_byteenable          (mm_interconnect_0_pixel_buffer_dma_avalon_control_slave_byteenable),          //                                               .byteenable
		.press_s1_address                                          (mm_interconnect_0_press_s1_address),                                          //                                       press_s1.address
		.press_s1_readdata                                         (mm_interconnect_0_press_s1_readdata),                                         //                                               .readdata
		.sdram_clk_pll_slave_address                               (mm_interconnect_0_sdram_clk_pll_slave_address),                               //                            sdram_clk_pll_slave.address
		.sdram_clk_pll_slave_write                                 (mm_interconnect_0_sdram_clk_pll_slave_write),                                 //                                               .write
		.sdram_clk_pll_slave_read                                  (mm_interconnect_0_sdram_clk_pll_slave_read),                                  //                                               .read
		.sdram_clk_pll_slave_readdata                              (mm_interconnect_0_sdram_clk_pll_slave_readdata),                              //                                               .readdata
		.sdram_clk_pll_slave_writedata                             (mm_interconnect_0_sdram_clk_pll_slave_writedata),                             //                                               .writedata
		.sdram_controller_0_s1_address                             (mm_interconnect_0_sdram_controller_0_s1_address),                             //                          sdram_controller_0_s1.address
		.sdram_controller_0_s1_write                               (mm_interconnect_0_sdram_controller_0_s1_write),                               //                                               .write
		.sdram_controller_0_s1_read                                (mm_interconnect_0_sdram_controller_0_s1_read),                                //                                               .read
		.sdram_controller_0_s1_readdata                            (mm_interconnect_0_sdram_controller_0_s1_readdata),                            //                                               .readdata
		.sdram_controller_0_s1_writedata                           (mm_interconnect_0_sdram_controller_0_s1_writedata),                           //                                               .writedata
		.sdram_controller_0_s1_byteenable                          (mm_interconnect_0_sdram_controller_0_s1_byteenable),                          //                                               .byteenable
		.sdram_controller_0_s1_readdatavalid                       (mm_interconnect_0_sdram_controller_0_s1_readdatavalid),                       //                                               .readdatavalid
		.sdram_controller_0_s1_waitrequest                         (mm_interconnect_0_sdram_controller_0_s1_waitrequest),                         //                                               .waitrequest
		.sdram_controller_0_s1_chipselect                          (mm_interconnect_0_sdram_controller_0_s1_chipselect)                           //                                               .chipselect
	);

	Video_System_irq_mapper irq_mapper (
		.clk        (clk_0),                              //       clk.clk
		.reset      (rst_controller_001_reset_out_reset), // clk_reset.reset
		.sender_irq (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_n),                       // reset_in0.reset
		.clk            (clk_0),                          //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_n),                               // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),      // reset_in1.reset
		.clk            (clk_0),                                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (video_pll_0_reset_source_reset),     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (video_pll_0_vga_clk_clk),            //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.reset_in1      (~reset_n),                           // reset_in1.reset
		.clk            (sdram_out_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
